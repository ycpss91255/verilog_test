module eazy_led (
  input  [9:0] iSW,
  output [9:0] oLED
);

assign oLED = iSW;

endmodule

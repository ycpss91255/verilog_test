module multiplexer (
  input [2:0] iClk,
  input [1:0] iSW,
  output      oClk
);



endmodule
